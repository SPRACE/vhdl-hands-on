-------------------------------------------------------------------------------
-- Title      : Patter Checker
-- Project    : 
-------------------------------------------------------------------------------
-- File       : pattern-checker.vhd
-- Author     : Vitor Finotti  <vfinotti@vfinotti-desktop.ncc.unesp.br>
-- Company    : Sao Paulo Research and Analysis Center,  SPRACE
-- Created    : 2018-02-08
-- Last update: 2018-02-08
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: In this this project, the LED will only blink when the push
-- buttons are pressed in a patter that matches the switches'.
-------------------------------------------------------------------------------
-- Copyright (c) 2018 Sao Paulo Research and Analysis Center,  SPRACE

-- This program is free software: you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public License
-- as published by the Free Software Foundation, either version 3 of
-- the License, or (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful, but
-- WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this program. If not, see
-- <http://www.gnu.org/licenses/>.
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2018-02-08  1.0      vfinotti        Created
-------------------------------------------------------------------------------

entity patter_checker_top is

    generic (
        g_input_width : natural := 3);  -- num of switches and push-buttons

    port (
        push_buttons_i : in  std_logic_vector(g_input_width-1 downto 0);
        switches_i     : in  std_logic_vector(g_input_width-1 downto 0);
        led_o          : out std_logic);

end entity patter_checker_top;

architecture rtl of pattern_checker_top is

begin  -- architecture rtl

    led_o <=     switches_i(0) and push_buttons_i(0)
             and switches_i(1) and push_buttons_i(1)
             and switches_i(2) and push_buttons_i(2);

end architecture rtl;
